-- SPI controller
  constant CFG_SPICTRL_ENABLE : integer := CONFIG_SPICTRL_ENABLE;

